// sort.v
//Lab 2 Part 4.2: Creating a Qsys component to sort

//Chris Bird, Lillie Deas, Kaila Balancio

module scroll (clock, resetn, KEY )
input clock;
input resetn;


always @ (posedge clock or posedge resetn)
begin
	if(resetn)

	else 
	begin


	end
end
endmodule
